library ieee;
use ieee.std_logic_1164.ALL;

entity top is
	port(
		-- PCIe #PERST
		pcie_nperst : in std_logic;

		-- PCIe refclk
		refclk : in std_logic;

		-- PCIe rx
		pcie_rx : in std_logic_vector(3 downto 0);

		-- PCIe tx
		pcie_tx : out std_logic_vector(3 downto 0);

		-- independent clock
		fixedclk_serdes : in std_logic
	);
end entity;

architecture rtl of top is
	-- async reset
	signal cpu_reset : std_logic;

	-- clock
	signal cpu_clk : std_logic;

	-- status
	signal cpu_halted : std_logic;

	-- instruction bus (Avalon-MM)
	signal cpu_i_addr : std_logic_vector(31 downto 0);
	signal cpu_i_rddata : std_logic_vector(63 downto 0);
	signal cpu_i_rdreq : std_logic;
	signal cpu_i_waitrequest : std_logic;

	-- data bus (Avalon-MM)
	signal cpu_d_addr : std_logic_vector(31 downto 0);
	signal cpu_d_rddata : std_logic_vector(31 downto 0);
	signal cpu_d_rdreq : std_logic;
	signal cpu_d_wrdata : std_logic_vector(31 downto 0);
	signal cpu_d_wrreq : std_logic;
	signal cpu_d_waitrequest : std_logic;

	component cpu is
		generic(
			address_width : integer
		);
		port(
			-- async reset
			reset : in std_logic;

			-- clock
			clk : in std_logic;

			-- status
			halted : out std_logic;

			-- instruction bus (Avalon-MM)
			i_addr : out std_logic_vector(31 downto 0);
			i_rddata : in std_logic_vector(63 downto 0);
			i_rdreq : out std_logic;
			i_waitrequest : in std_logic;

			-- data bus (Avalon-MM)
			d_addr : out std_logic_vector(31 downto 0);
			d_rddata : in std_logic_vector(31 downto 0);
			d_rdreq : out std_logic;
			d_wrdata : out std_logic_vector(31 downto 0);
			d_wrreq : out std_logic;
			d_waitrequest : in std_logic
		);
	end component;

	-- clocks
	signal pld_clk : std_logic;
	signal core_clk_out : std_logic;
	signal cal_blk_clk : std_logic;

	signal app_clk : std_logic;			-- application clock

	-- PCIe internal rx interface (Avalon-ST), synchronous to app_clk
	signal pcie_rx_ready : std_logic;
	signal pcie_rx_valid : std_logic;
	signal pcie_rx_data : std_logic_vector(63 downto 0);
	signal pcie_rx_sop : std_logic;
	signal pcie_rx_eop : std_logic;
	signal pcie_rx_err : std_logic;

	signal pcie_rx_mask : std_logic;
	signal pcie_rx_bardec : std_logic_vector(7 downto 0);

	-- PCIe internal tx interface (Avalon-ST), synchronous to app_clk
	signal pcie_tx_ready : std_logic;
	signal pcie_tx_valid : std_logic;
	signal pcie_tx_data : std_logic_vector(63 downto 0);
	signal pcie_tx_sop : std_logic;
	signal pcie_tx_eop : std_logic;
	signal pcie_tx_err : std_logic;

	-- completion interface
	signal cpl_pending : std_logic;

	-- interrupts
	signal app_int_sts : std_logic;
	signal app_int_ack : std_logic;

	signal app_msi_req : std_logic;
	signal app_msi_num : std_logic_vector(4 downto 0);
	signal app_msi_tc : std_logic_vector(2 downto 0);
	signal app_msi_ack : std_logic;

	-- reset
	signal npor : std_logic;	-- power on reset (external)
	signal app_rstn : std_logic;	-- application reset (generated by reset controller)
	signal srst : std_logic;	-- datapath reset (generated by reset controller)
	signal crst : std_logic;	-- configuration space reset (generated by reset controller)

	-- transceiver state
	signal dlup_exit : std_logic;
	signal hotrst_exit : std_logic;
	signal l2_exit : std_logic;
	signal ltssm : std_logic_vector(4 downto 0);
	signal rc_pll_locked : std_logic;
	signal reset_status : std_logic;
	signal suc_spd_neg : std_logic;

	-- PHY reconfiguration interface
	signal reconfig_clk : std_logic;
	signal reconfig_busy : std_logic;
	signal reconfig_fromgxb : std_logic_vector(4 downto 0);
	signal reconfig_togxb : std_logic_vector(3 downto 0);

	-- power management
	signal gxb_powerdown : std_logic;
	signal pll_powerdown : std_logic;
	signal pm_auxpwr : std_logic;
	signal pm_data : std_logic_vector(9 downto 0);
	signal pm_event : std_logic;
	signal pme_to_cr : std_logic;
	signal pme_to_sr : std_logic;

	-- local management interface
	signal lmi_addr : std_logic_vector(11 downto 0);
	signal lmi_rden : std_logic;
	signal lmi_din : std_logic_vector(31 downto 0);
	signal lmi_wren : std_logic;
	signal lmi_dout : std_logic_vector(31 downto 0);
	signal lmi_ack : std_logic;

	-- configuration space
	signal tl_cfg_add : std_logic_vector(3 downto 0);
	signal tl_cfg_ctl : std_logic_vector(31 downto 0);
	signal tl_cfg_ctl_wr : std_logic;
	signal tl_cfg_sts : std_logic_vector(52 downto 0);
	signal tl_cfg_sts_wr : std_logic;
begin
	cpu_reset <= '1';
	cpu_clk <= '0';

	cpu_i_rddata <= (others => '0');
	cpu_i_waitrequest <= '1';

	cpu_d_rddata <= (others => '0');
	cpu_d_waitrequest <= '1';

	c : cpu
		generic map(
			address_width => 32
		)
		port map(
			reset => cpu_reset,
			clk => cpu_clk,
			halted => cpu_halted,
			i_addr => cpu_i_addr,
			i_rddata => cpu_i_rddata,
			i_rdreq => cpu_i_rdreq,
			i_waitrequest => cpu_i_waitrequest,
			d_addr => cpu_d_addr,
			d_rddata => cpu_d_rddata,
			d_rdreq => cpu_d_rdreq,
			d_wrdata => cpu_d_wrdata,
			d_wrreq => cpu_d_wrreq,
			d_waitrequest => cpu_d_waitrequest
		);

	-- clocks
	pld_clk <= core_clk_out;		-- needs to be connected
	app_clk <= pld_clk;			-- app is synchronous to pld_clk
	cal_blk_clk <= core_clk_out;

	-- PCIe internal rx interface (Avalon-ST)
	pcie_rx_ready <= '0';
	pcie_rx_mask <= '0';

	-- PCIe internal tx interface (Avalon-ST)
	pcie_tx_valid <= '0';
	pcie_tx_data <= (others => '0');
	pcie_tx_sop <= '0';
	pcie_tx_eop <= '0';
	pcie_tx_err <= '0';

	-- completion interface
	cpl_pending <= '0';

	-- interrupts
	app_int_sts <= '0';

	app_msi_req <= '0';
	app_msi_num <= (others => '0');
	app_msi_tc <= (others => '0');

	-- reset
	npor <= pcie_nperst;

	-- power management
	gxb_powerdown <= '0';
	pll_powerdown <= '0';
	pm_auxpwr <= '0';
	pm_data <= (others => '0');		-- todo
	pm_event <= '0';
	pme_to_cr <= '0';

	-- local management interface
	lmi_addr <= (others => '0');
	lmi_rden <= '0';
	lmi_din <= (others => '0');
	lmi_wren <= '0';

	pcie_inst : entity work.pcie
		port map (
			-- external PCIe interface
			rx_in0 => pcie_rx(0),
			rx_in1 => pcie_rx(1),
			rx_in2 => pcie_rx(2),
			rx_in3 => pcie_rx(3),
			tx_out0 => pcie_tx(0),
			tx_out1 => pcie_tx(1),
			tx_out2 => pcie_tx(2),
			tx_out3 => pcie_tx(3),

			-- clocks
			refclk => refclk,
			fixedclk_serdes => fixedclk_serdes,
			pclk_in => '0',				-- PIPE simulation only
			pld_clk => pld_clk,
			core_clk_out => core_clk_out,

			-- PCIe internal rx interface (Avalon-ST)
			rx_st_ready0 => pcie_rx_ready,
			rx_st_valid0 => pcie_rx_valid,
			rx_st_data0 => pcie_rx_data,
			rx_st_sop0 => pcie_rx_sop,
			rx_st_eop0 => pcie_rx_eop,
			rx_st_err0 => pcie_rx_err,

			rx_st_mask0 => pcie_rx_mask,
			rx_st_bardec0 => pcie_rx_bardec,
			rx_st_be0 => open,			-- deprecated

			-- PCIe internal tx interface (Avalon-ST)
			tx_st_ready0 => pcie_tx_ready,
			tx_st_valid0 => pcie_tx_valid,
			tx_st_data0 => pcie_tx_data,
			tx_st_sop0 => pcie_tx_sop,
			tx_st_eop0 => pcie_tx_eop,
			tx_st_err0 => pcie_tx_err,

			-- completion interface
			cpl_err => (others => '0'),		-- todo
			cpl_pending => cpl_pending,
			ko_cpl_spc_vc0 => open,			-- todo

			-- interrupts
			app_int_sts => app_int_sts,
			app_int_ack => app_int_ack,
			app_msi_req => app_msi_req,
			app_msi_num => app_msi_num,
			app_msi_tc => app_msi_tc,
			app_msi_ack => app_msi_ack,
			pex_msi_num => (others => '0'),		-- todo

			-- reset
			npor => npor,
			crst => crst,
			srst => srst,

			-- transceiver state
			dlup_exit => dlup_exit,
			hotrst_exit => hotrst_exit,
			l2_exit => l2_exit,
			ltssm => ltssm,
			rc_pll_locked => rc_pll_locked,
			reset_status => reset_status,
			suc_spd_neg => suc_spd_neg,
			rc_rx_digitalreset => open,

			-- PHY reconfiguration interface
			busy_altgxb_reconfig => reconfig_busy,
			cal_blk_clk => cal_blk_clk,
			reconfig_clk => reconfig_clk,
			reconfig_togxb => reconfig_togxb,
			reconfig_fromgxb => reconfig_fromgxb,

			-- power management
			gxb_powerdown => gxb_powerdown,
			pll_powerdown => pll_powerdown,
			pm_auxpwr => pm_auxpwr,
			pm_data => pm_data,
			pm_event => pm_event,
			pme_to_cr => pme_to_cr,
			pme_to_sr => pme_to_sr,

			-- local management interface
			lmi_addr => lmi_addr,
			lmi_din => lmi_din,
			lmi_rden => lmi_rden,
			lmi_wren => lmi_wren,
			lmi_ack => lmi_ack,
			lmi_dout => lmi_dout,

			-- configuration space
			tl_cfg_add => tl_cfg_add,
			tl_cfg_ctl => tl_cfg_ctl,
			tl_cfg_ctl_wr => tl_cfg_ctl_wr,
			tl_cfg_sts => tl_cfg_sts,
			tl_cfg_sts_wr => tl_cfg_sts_wr,

			-- PCIe credits (todo)
			tx_cred0 => open,

			-- ECC error handling (todo)
			derr_cor_ext_rcv0 => open,
			derr_cor_ext_rpl => open,
			derr_rpl => open,
			r2c_err0 => open,

			-- test interface (unused)
			test_in => (others => '0'),
			lane_act => open,

			-- simulation only (do not work on actual hardware)
			clk250_out => open,
			clk500_out => open,

			-- debug signals
			rx_fifo_empty0 => open,
			rx_fifo_full0 => open,
			tx_fifo_empty0 => open,
			tx_fifo_full0 => open,
			tx_fifo_rdptr0 => open,
			tx_fifo_wrptr0 => open,

			-- PIPE mode (disabled)
			pipe_mode => '0',

			hpg_ctrler => (others => '0'),
			phystatus_ext => '0',
			rxdata0_ext => (others => '0'),
			rxdata1_ext => (others => '0'),
			rxdata2_ext => (others => '0'),
			rxdata3_ext => (others => '0'),
			rxdatak0_ext => '0',
			rxdatak1_ext => '0',
			rxdatak2_ext => '0',
			rxdatak3_ext => '0',
			rxelecidle0_ext => '0',
			rxelecidle1_ext => '0',
			rxelecidle2_ext => '0',
			rxelecidle3_ext => '0',
			rxstatus0_ext => (others => '0'),
			rxstatus1_ext => (others => '0'),
			rxstatus2_ext => (others => '0'),
			rxstatus3_ext => (others => '0'),
			rxvalid0_ext => '0',
			rxvalid1_ext => '0',
			rxvalid2_ext => '0',
			rxvalid3_ext => '0',

			rate_ext => open,
			rxpolarity0_ext => open,
			rxpolarity1_ext => open,
			rxpolarity2_ext => open,
			rxpolarity3_ext => open,
			txcompl0_ext => open,
			txcompl1_ext => open,
			txcompl2_ext => open,
			txcompl3_ext => open,
			txdata0_ext => open,
			txdata1_ext => open,
			txdata2_ext => open,
			txdata3_ext => open,
			txdatak0_ext => open,
			txdatak1_ext => open,
			txdatak2_ext => open,
			txdatak3_ext => open,
			txdetectrx_ext => open,
			txelecidle0_ext => open,
			txelecidle1_ext => open,
			txelecidle2_ext => open,
			txelecidle3_ext => open
		);

	pll_inst : entity work.pll
		port map (
			inclk0 => fixedclk_serdes,
			c0 => reconfig_clk
		);

	pcie_reset_inst : entity work.pcie_rs_hip
		port map (
			-- power on reset (external, low active)
			npor => npor,

			-- clock
			pld_clk => pld_clk,

			-- current transceiver state
			dlup_exit => dlup_exit,		-- data link up
			hotrst_exit => hotrst_exit,	-- hot reset
			l2_exit => l2_exit,		-- layer 2
			ltssm => ltssm,			-- link training state machine

			-- generated reset signals
			app_rstn => app_rstn,		-- generated app reset (low active)
			crst => crst,			-- generated crst
			srst => srst,			-- generated srst

			test_sim => '0'
		);

	pcie_reconfig_inst : entity work.pcie_reconfig
		port map (
			reconfig_clk => reconfig_clk,
			busy => reconfig_busy,
			reconfig_fromgxb => reconfig_fromgxb,
			reconfig_togxb => reconfig_togxb
		);
end architecture;

library work;
use work.ALL;

configuration rtl of top is
	for rtl
		for c : cpu
			use entity work.cpu_sequential;
			for rtl
				for register_file : registers
					use entity work.altera_registers;
				end for;
			end for;
		end for;
	end for;
end configuration;
