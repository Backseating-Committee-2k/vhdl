-- megafunction wizard: %ALTGX%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: alt_c3gxb 

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV GX"
-- Retrieval info: PRIVATE: IP_MODE STRING "PCIE_HIP_8"
-- Retrieval info: PRIVATE: LOCKDOWN_EXCL STRING "PCIE"
-- Retrieval info: PRIVATE: NUM_KEYS NUMERIC "0"
-- Retrieval info: PRIVATE: RECONFIG_PROTOCOL STRING "BASIC"
-- Retrieval info: PRIVATE: RECONFIG_SUBPROTOCOL STRING "none"
-- Retrieval info: PRIVATE: RX_ENABLE_DC_COUPLING STRING "false"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: WIZ_BASE_DATA_RATE STRING "2500"
-- Retrieval info: PRIVATE: WIZ_BASE_DATA_RATE_ENABLE STRING "0"
-- Retrieval info: PRIVATE: WIZ_DATA_RATE STRING "2500"
-- Retrieval info: PRIVATE: WIZ_DPRIO_INCLK_FREQ_ARRAY STRING "100 100 100 100 100 100 100 100 100 100 100 100 100 100 100 100 100 100 100 100"
-- Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_A STRING "2000"
-- Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_A_UNIT STRING "Mbps"
-- Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_B STRING "100"
-- Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_B_UNIT STRING "MHz"
-- Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_SELECTION NUMERIC "0"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK0_FREQ STRING "100.0"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK0_PROTOCOL STRING "PCI Express (PIPE)"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK1_FREQ STRING "250"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK1_PROTOCOL STRING "Basic"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK2_FREQ STRING "250"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK2_PROTOCOL STRING "Basic"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK3_FREQ STRING "250"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK3_PROTOCOL STRING "Basic"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK4_FREQ STRING "250"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK4_PROTOCOL STRING "Basic"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK5_FREQ STRING "250"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK5_PROTOCOL STRING "Basic"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK6_FREQ STRING "250"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK6_PROTOCOL STRING "Basic"
-- Retrieval info: PRIVATE: WIZ_ENABLE_EQUALIZER_CTRL NUMERIC "1"
-- Retrieval info: PRIVATE: WIZ_EQUALIZER_CTRL_SETTING NUMERIC "1"
-- Retrieval info: PRIVATE: WIZ_FORCE_DEFAULT_SETTINGS NUMERIC "0"
-- Retrieval info: PRIVATE: WIZ_INCLK_FREQ STRING "100.0"
-- Retrieval info: PRIVATE: WIZ_INCLK_FREQ_ARRAY STRING "100.0 125.0"
-- Retrieval info: PRIVATE: WIZ_INPUT_A STRING "2500"
-- Retrieval info: PRIVATE: WIZ_INPUT_A_UNIT STRING "Mbps"
-- Retrieval info: PRIVATE: WIZ_INPUT_B STRING "100.0"
-- Retrieval info: PRIVATE: WIZ_INPUT_B_UNIT STRING "MHz"
-- Retrieval info: PRIVATE: WIZ_INPUT_SELECTION NUMERIC "0"
-- Retrieval info: PRIVATE: WIZ_PROTOCOL STRING "PCI Express (PIPE)"
-- Retrieval info: PRIVATE: WIZ_SUBPROTOCOL STRING "Gen 1-x4"
-- Retrieval info: PRIVATE: WIZ_WORD_ALIGN_FLIP_PATTERN STRING "0"
-- Retrieval info: PARAMETER: STARTING_CHANNEL_NUMBER NUMERIC "0"
-- Retrieval info: CONSTANT: EFFECTIVE_DATA_RATE STRING "2500 Mbps"
-- Retrieval info: CONSTANT: ENABLE_LC_TX_PLL STRING "false"
-- Retrieval info: CONSTANT: ENABLE_PLL_INCLK_ALT_DRIVE_RX_CRU STRING "true"
-- Retrieval info: CONSTANT: ENABLE_PLL_INCLK_DRIVE_RX_CRU STRING "true"
-- Retrieval info: CONSTANT: EQUALIZER_DCGAIN_SETTING NUMERIC "1"
-- Retrieval info: CONSTANT: GEN_RECONFIG_PLL STRING "false"
-- Retrieval info: CONSTANT: GX_CHANNEL_TYPE STRING ""
-- Retrieval info: CONSTANT: INPUT_CLOCK_FREQUENCY STRING "100.0 MHz"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone IV GX"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_SPEED_GRADE STRING "6"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_VARIANT STRING "ANY"
-- Retrieval info: CONSTANT: LOOPBACK_MODE STRING "none"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "alt_c3gxb"
-- Retrieval info: CONSTANT: NUMBER_OF_CHANNELS NUMERIC "4"
-- Retrieval info: CONSTANT: OPERATION_MODE STRING "duplex"
-- Retrieval info: CONSTANT: PLL_BANDWIDTH_TYPE STRING "Auto"
-- Retrieval info: CONSTANT: PLL_CONTROL_WIDTH NUMERIC "1"
-- Retrieval info: CONSTANT: PLL_INCLK_PERIOD NUMERIC "10000"
-- Retrieval info: CONSTANT: PLL_PFD_FB_MODE STRING "internal"
-- Retrieval info: CONSTANT: PREEMPHASIS_CTRL_1STPOSTTAP_SETTING NUMERIC "1"
-- Retrieval info: CONSTANT: PROTOCOL STRING "pcie"
-- Retrieval info: CONSTANT: RECEIVER_TERMINATION STRING "oct_100_ohms"
-- Retrieval info: CONSTANT: RECONFIG_DPRIO_MODE NUMERIC "0"
-- Retrieval info: CONSTANT: RX_8B_10B_MODE STRING "normal"
-- Retrieval info: CONSTANT: RX_ALIGN_PATTERN STRING "0101111100"
-- Retrieval info: CONSTANT: RX_ALIGN_PATTERN_LENGTH NUMERIC "10"
-- Retrieval info: CONSTANT: RX_ALLOW_ALIGN_POLARITY_INVERSION STRING "false"
-- Retrieval info: CONSTANT: RX_ALLOW_PIPE_POLARITY_INVERSION STRING "true"
-- Retrieval info: CONSTANT: RX_BITSLIP_ENABLE STRING "false"
-- Retrieval info: CONSTANT: RX_BYTE_ORDERING_MODE STRING "NONE"
-- Retrieval info: CONSTANT: RX_CHANNEL_BONDING STRING "x4"
-- Retrieval info: CONSTANT: RX_CHANNEL_WIDTH NUMERIC "8"
-- Retrieval info: CONSTANT: RX_COMMON_MODE STRING "0.82v"
-- Retrieval info: CONSTANT: RX_CRU_INCLOCK0_PERIOD NUMERIC "10000"
-- Retrieval info: CONSTANT: RX_DATAPATH_PROTOCOL STRING "pipe"
-- Retrieval info: CONSTANT: RX_DATA_RATE NUMERIC "2500"
-- Retrieval info: CONSTANT: RX_DATA_RATE_REMAINDER NUMERIC "0"
-- Retrieval info: CONSTANT: RX_DIGITALRESET_PORT_WIDTH NUMERIC "1"
-- Retrieval info: CONSTANT: RX_ENABLE_BIT_REVERSAL STRING "false"
-- Retrieval info: CONSTANT: RX_ENABLE_LOCK_TO_DATA_SIG STRING "false"
-- Retrieval info: CONSTANT: RX_ENABLE_LOCK_TO_REFCLK_SIG STRING "false"
-- Retrieval info: CONSTANT: RX_ENABLE_SELF_TEST_MODE STRING "false"
-- Retrieval info: CONSTANT: RX_FORCE_SIGNAL_DETECT STRING "false"
-- Retrieval info: CONSTANT: RX_PPMSELECT NUMERIC "8"
-- Retrieval info: CONSTANT: RX_RATE_MATCH_FIFO_MODE STRING "normal"
-- Retrieval info: CONSTANT: RX_RATE_MATCH_PATTERN1 STRING "11010000111010000011"
-- Retrieval info: CONSTANT: RX_RATE_MATCH_PATTERN2 STRING "00101111000101111100"
-- Retrieval info: CONSTANT: RX_RATE_MATCH_PATTERN_SIZE NUMERIC "20"
-- Retrieval info: CONSTANT: RX_RUN_LENGTH NUMERIC "40"
-- Retrieval info: CONSTANT: RX_RUN_LENGTH_ENABLE STRING "true"
-- Retrieval info: CONSTANT: RX_SIGNAL_DETECT_THRESHOLD NUMERIC "4"
-- Retrieval info: CONSTANT: RX_USE_ALIGN_STATE_MACHINE STRING "true"
-- Retrieval info: CONSTANT: RX_USE_CLKOUT STRING "false"
-- Retrieval info: CONSTANT: RX_USE_CORECLK STRING "false"
-- Retrieval info: CONSTANT: RX_USE_DESERIALIZER_DOUBLE_DATA_MODE STRING "false"
-- Retrieval info: CONSTANT: RX_USE_DESKEW_FIFO STRING "false"
-- Retrieval info: CONSTANT: RX_USE_DOUBLE_DATA_MODE STRING "false"
-- Retrieval info: CONSTANT: RX_USE_PIPE8B10BINVPOLARITY STRING "true"
-- Retrieval info: CONSTANT: RX_USE_RATE_MATCH_PATTERN1_ONLY STRING "false"
-- Retrieval info: CONSTANT: TRANSMITTER_TERMINATION STRING "oct_100_ohms"
-- Retrieval info: CONSTANT: TX_8B_10B_MODE STRING "normal"
-- Retrieval info: CONSTANT: TX_ALLOW_POLARITY_INVERSION STRING "false"
-- Retrieval info: CONSTANT: TX_CHANNEL_BONDING STRING "x4"
-- Retrieval info: CONSTANT: TX_CHANNEL_WIDTH NUMERIC "8"
-- Retrieval info: CONSTANT: TX_CLKOUT_WIDTH NUMERIC "4"
-- Retrieval info: CONSTANT: TX_COMMON_MODE STRING "0.65v"
-- Retrieval info: CONSTANT: TX_DATA_RATE NUMERIC "2500"
-- Retrieval info: CONSTANT: TX_DATA_RATE_REMAINDER NUMERIC "0"
-- Retrieval info: CONSTANT: TX_DIGITALRESET_PORT_WIDTH NUMERIC "1"
-- Retrieval info: CONSTANT: TX_ENABLE_BIT_REVERSAL STRING "false"
-- Retrieval info: CONSTANT: TX_ENABLE_SELF_TEST_MODE STRING "false"
-- Retrieval info: CONSTANT: TX_PLL_BANDWIDTH_TYPE STRING "Auto"
-- Retrieval info: CONSTANT: TX_PLL_INCLK0_PERIOD NUMERIC "10000"
-- Retrieval info: CONSTANT: TX_PLL_TYPE STRING "CMU"
-- Retrieval info: CONSTANT: TX_SLEW_RATE STRING "low"
-- Retrieval info: CONSTANT: TX_TRANSMIT_PROTOCOL STRING "pipe"
-- Retrieval info: CONSTANT: TX_USE_CORECLK STRING "false"
-- Retrieval info: CONSTANT: TX_USE_DOUBLE_DATA_MODE STRING "false"
-- Retrieval info: CONSTANT: TX_USE_SERIALIZER_DOUBLE_DATA_MODE STRING "false"
-- Retrieval info: CONSTANT: USE_CALIBRATION_BLOCK STRING "true"
-- Retrieval info: CONSTANT: VOD_CTRL_SETTING NUMERIC "4"
-- Retrieval info: CONSTANT: coreclkout_control_width NUMERIC "1"
-- Retrieval info: CONSTANT: elec_idle_infer_enable STRING "false"
-- Retrieval info: CONSTANT: enable_0ppm STRING "false"
-- Retrieval info: CONSTANT: equalization_setting NUMERIC "5"
-- Retrieval info: CONSTANT: gxb_powerdown_width NUMERIC "1"
-- Retrieval info: CONSTANT: hip_enable STRING "true"
-- Retrieval info: CONSTANT: iqtxrxclk_allowed STRING ""
-- Retrieval info: CONSTANT: number_of_quads NUMERIC "1"
-- Retrieval info: CONSTANT: pll_divide_by STRING "2"
-- Retrieval info: CONSTANT: pll_multiply_by STRING "25"
-- Retrieval info: CONSTANT: reconfig_calibration STRING "true"
-- Retrieval info: CONSTANT: reconfig_fromgxb_port_width NUMERIC "5"
-- Retrieval info: CONSTANT: reconfig_pll_control_width NUMERIC "1"
-- Retrieval info: CONSTANT: reconfig_togxb_port_width NUMERIC "4"
-- Retrieval info: CONSTANT: rx_cdrctrl_enable STRING "true"
-- Retrieval info: CONSTANT: rx_deskew_pattern STRING "0"
-- Retrieval info: CONSTANT: rx_dwidth_factor NUMERIC "1"
-- Retrieval info: CONSTANT: rx_enable_second_order_loop STRING "false"
-- Retrieval info: CONSTANT: rx_loop_1_digital_filter NUMERIC "8"
-- Retrieval info: CONSTANT: rx_signal_detect_loss_threshold STRING "3"
-- Retrieval info: CONSTANT: rx_signal_detect_valid_threshold STRING "14"
-- Retrieval info: CONSTANT: rx_use_external_termination STRING "false"
-- Retrieval info: CONSTANT: rx_word_aligner_num_byte NUMERIC "1"
-- Retrieval info: CONSTANT: top_module_name STRING "pcie_serdes"
-- Retrieval info: CONSTANT: tx_bitslip_enable STRING "FALSE"
-- Retrieval info: CONSTANT: tx_dwidth_factor NUMERIC "1"
-- Retrieval info: CONSTANT: tx_use_external_termination STRING "false"
-- Retrieval info: USED_PORT: cal_blk_clk 0 0 0 0 INPUT NODEFVAL "cal_blk_clk"
-- Retrieval info: USED_PORT: coreclkout 0 0 1 0 OUTPUT NODEFVAL "coreclkout[0..0]"
-- Retrieval info: USED_PORT: fixedclk 0 0 0 0 INPUT NODEFVAL "fixedclk"
-- Retrieval info: USED_PORT: gxb_powerdown 0 0 1 0 INPUT NODEFVAL "gxb_powerdown[0..0]"
-- Retrieval info: USED_PORT: hip_tx_clkout 0 0 4 0 OUTPUT NODEFVAL "hip_tx_clkout[3..0]"
-- Retrieval info: USED_PORT: pipe8b10binvpolarity 0 0 4 0 INPUT NODEFVAL "pipe8b10binvpolarity[3..0]"
-- Retrieval info: USED_PORT: pipedatavalid 0 0 4 0 OUTPUT NODEFVAL "pipedatavalid[3..0]"
-- Retrieval info: USED_PORT: pipeelecidle 0 0 4 0 OUTPUT NODEFVAL "pipeelecidle[3..0]"
-- Retrieval info: USED_PORT: pipephydonestatus 0 0 4 0 OUTPUT NODEFVAL "pipephydonestatus[3..0]"
-- Retrieval info: USED_PORT: pipestatus 0 0 12 0 OUTPUT NODEFVAL "pipestatus[11..0]"
-- Retrieval info: USED_PORT: pll_areset 0 0 1 0 INPUT NODEFVAL "pll_areset[0..0]"
-- Retrieval info: USED_PORT: pll_inclk 0 0 1 0 INPUT NODEFVAL "pll_inclk[0..0]"
-- Retrieval info: USED_PORT: pll_locked 0 0 1 0 OUTPUT NODEFVAL "pll_locked[0..0]"
-- Retrieval info: USED_PORT: powerdn 0 0 8 0 INPUT NODEFVAL "powerdn[7..0]"
-- Retrieval info: USED_PORT: reconfig_clk 0 0 0 0 INPUT NODEFVAL "reconfig_clk"
-- Retrieval info: USED_PORT: reconfig_fromgxb 0 0 5 0 OUTPUT NODEFVAL "reconfig_fromgxb[4..0]"
-- Retrieval info: USED_PORT: reconfig_togxb 0 0 4 0 INPUT NODEFVAL "reconfig_togxb[3..0]"
-- Retrieval info: USED_PORT: rx_analogreset 0 0 1 0 INPUT NODEFVAL "rx_analogreset[0..0]"
-- Retrieval info: USED_PORT: rx_ctrldetect 0 0 4 0 OUTPUT NODEFVAL "rx_ctrldetect[3..0]"
-- Retrieval info: USED_PORT: rx_datain 0 0 4 0 INPUT NODEFVAL "rx_datain[3..0]"
-- Retrieval info: USED_PORT: rx_dataout 0 0 32 0 OUTPUT NODEFVAL "rx_dataout[31..0]"
-- Retrieval info: USED_PORT: rx_digitalreset 0 0 1 0 INPUT NODEFVAL "rx_digitalreset[0..0]"
-- Retrieval info: USED_PORT: rx_elecidleinfersel 0 0 12 0 INPUT NODEFVAL "rx_elecidleinfersel[11..0]"
-- Retrieval info: USED_PORT: rx_freqlocked 0 0 4 0 OUTPUT NODEFVAL "rx_freqlocked[3..0]"
-- Retrieval info: USED_PORT: rx_patterndetect 0 0 4 0 OUTPUT NODEFVAL "rx_patterndetect[3..0]"
-- Retrieval info: USED_PORT: rx_syncstatus 0 0 4 0 OUTPUT NODEFVAL "rx_syncstatus[3..0]"
-- Retrieval info: USED_PORT: tx_ctrlenable 0 0 4 0 INPUT NODEFVAL "tx_ctrlenable[3..0]"
-- Retrieval info: USED_PORT: tx_datain 0 0 32 0 INPUT NODEFVAL "tx_datain[31..0]"
-- Retrieval info: USED_PORT: tx_dataout 0 0 4 0 OUTPUT NODEFVAL "tx_dataout[3..0]"
-- Retrieval info: USED_PORT: tx_detectrxloop 0 0 4 0 INPUT NODEFVAL "tx_detectrxloop[3..0]"
-- Retrieval info: USED_PORT: tx_digitalreset 0 0 1 0 INPUT NODEFVAL "tx_digitalreset[0..0]"
-- Retrieval info: USED_PORT: tx_forcedispcompliance 0 0 4 0 INPUT NODEFVAL "tx_forcedispcompliance[3..0]"
-- Retrieval info: USED_PORT: tx_forceelecidle 0 0 4 0 INPUT NODEFVAL "tx_forceelecidle[3..0]"
-- Retrieval info: CONNECT: @cal_blk_clk 0 0 0 0 cal_blk_clk 0 0 0 0
-- Retrieval info: CONNECT: @fixedclk 0 0 0 0 fixedclk 0 0 0 0
-- Retrieval info: CONNECT: @gxb_powerdown 0 0 1 0 gxb_powerdown 0 0 1 0
-- Retrieval info: CONNECT: @pipe8b10binvpolarity 0 0 4 0 pipe8b10binvpolarity 0 0 4 0
-- Retrieval info: CONNECT: @pll_areset 0 0 1 0 pll_areset 0 0 1 0
-- Retrieval info: CONNECT: @pll_inclk 0 0 1 0 pll_inclk 0 0 1 0
-- Retrieval info: CONNECT: @powerdn 0 0 8 0 powerdn 0 0 8 0
-- Retrieval info: CONNECT: @reconfig_clk 0 0 0 0 reconfig_clk 0 0 0 0
-- Retrieval info: CONNECT: @reconfig_togxb 0 0 4 0 reconfig_togxb 0 0 4 0
-- Retrieval info: CONNECT: @rx_analogreset 0 0 1 0 rx_analogreset 0 0 1 0
-- Retrieval info: CONNECT: @rx_datain 0 0 4 0 rx_datain 0 0 4 0
-- Retrieval info: CONNECT: @rx_digitalreset 0 0 1 0 rx_digitalreset 0 0 1 0
-- Retrieval info: CONNECT: @rx_elecidleinfersel 0 0 12 0 rx_elecidleinfersel 0 0 12 0
-- Retrieval info: CONNECT: @tx_ctrlenable 0 0 4 0 tx_ctrlenable 0 0 4 0
-- Retrieval info: CONNECT: @tx_datain 0 0 32 0 tx_datain 0 0 32 0
-- Retrieval info: CONNECT: @tx_detectrxloop 0 0 4 0 tx_detectrxloop 0 0 4 0
-- Retrieval info: CONNECT: @tx_digitalreset 0 0 1 0 tx_digitalreset 0 0 1 0
-- Retrieval info: CONNECT: @tx_forcedispcompliance 0 0 4 0 tx_forcedispcompliance 0 0 4 0
-- Retrieval info: CONNECT: @tx_forceelecidle 0 0 4 0 tx_forceelecidle 0 0 4 0
-- Retrieval info: CONNECT: coreclkout 0 0 1 0 @coreclkout 0 0 1 0
-- Retrieval info: CONNECT: hip_tx_clkout 0 0 4 0 @hip_tx_clkout 0 0 4 0
-- Retrieval info: CONNECT: pipedatavalid 0 0 4 0 @pipedatavalid 0 0 4 0
-- Retrieval info: CONNECT: pipeelecidle 0 0 4 0 @pipeelecidle 0 0 4 0
-- Retrieval info: CONNECT: pipephydonestatus 0 0 4 0 @pipephydonestatus 0 0 4 0
-- Retrieval info: CONNECT: pipestatus 0 0 12 0 @pipestatus 0 0 12 0
-- Retrieval info: CONNECT: pll_locked 0 0 1 0 @pll_locked 0 0 1 0
-- Retrieval info: CONNECT: reconfig_fromgxb 0 0 5 0 @reconfig_fromgxb 0 0 5 0
-- Retrieval info: CONNECT: rx_ctrldetect 0 0 4 0 @rx_ctrldetect 0 0 4 0
-- Retrieval info: CONNECT: rx_dataout 0 0 32 0 @rx_dataout 0 0 32 0
-- Retrieval info: CONNECT: rx_freqlocked 0 0 4 0 @rx_freqlocked 0 0 4 0
-- Retrieval info: CONNECT: rx_patterndetect 0 0 4 0 @rx_patterndetect 0 0 4 0
-- Retrieval info: CONNECT: rx_syncstatus 0 0 4 0 @rx_syncstatus 0 0 4 0
-- Retrieval info: CONNECT: tx_dataout 0 0 4 0 @tx_dataout 0 0 4 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL pcie_serdes.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL pcie_serdes.ppf TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL pcie_serdes.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL pcie_serdes.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL pcie_serdes.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL pcie_serdes_inst.vhd FALSE
